`include "dispatch_if.vh"
`include "types_pkg.vh"

module dispatch(
    input logic CLK, nRST,
    dispatch_if.DI diif
);

    import types_pkg::*;

    dispatch_t n_dispatch;
    dispatch_t dispatch;

    // hazards
    logic WAW_h;
    logic struct_h;
    logic hazard;

    logic [31:0] Instruction;
    opcode_t op;
    logic [4:0] rs, rt, rd;
    logic [15:0] imm;

    always_ff @ (posedge CLK, negedge nRST) begin: Pipeline_Latching
      if (~nRST)
        diif.out <= '0;
    	else
        diif.out <= n_dispatch;
    end

    always_comb begin : Pipeline_Output
      case (1'b1)
        diif.flush:  n_dispatch = '0;
        diif.freeze: n_dispatch = diif.out;
        hazard:      n_dispatch = diif.out;
        diif.ihit:   n_dispatch = dispatch;
        default:     n_dispatch = diif.out;
      endcase
    end

    always_comb begin: Instruction_Signals
      Instruction = diif.fetch.imemload;
      op = opcode_t'(Instruction[31:26]);
      rs = Instruction[25:21];
      rt = Instruction[20:16];
      rd = Instruction[15:11];
      imm = Instruction[15:0];
      func = funct_t'(Instruction[5:0]);
    end

    always_comb begin : Hazard_Logic
      case (cuif.cu.fu)
        ALU: struct_h = fust.alu.busy;
        LDST: struct_h = fust.ldst.busy;
        BRANCH: struct_h = fust.branch.busy;
        default: struct_h = 1'b0;
      endcase
      WAW_h = rst[rd].busy;
      hazard = struct_h | WAW_h;
    end

    always_comb begin : Dispatch_Out
      dispatch = diif.fetch.out;
      dispatch.hazard = hazard;
      dispatch.cu = cuif.cu;
    end

endmodule
