`ifndef DISPATCH_IF_VH
`define DISPATCH_IF_VH
`include "datapath_types.vh"

interface dispatch_if;
    import datapath_pkg::*;

    //Inputs from fetch
    typedef logic [2:0] fetch_t;
    fetch_t fetch;

    // Inputs to latch
    logic flush, freeze;

    // Inputs from issue 
    fust_s_t fust_s;
    fust_m_t fust_m;
    fust_g_t fust_g;

    // Inputs from writeback
    wb_t wb;
    
    // Inputs from memory
    logic ihit;
    
    // Outputs of stage
    dispatch_t out;
    
    modport DI (
        input fetch, flush, freeze, fust_s, fust_m, fust_g, wb, ihit,
        output out
    );

endinterface
`endif
