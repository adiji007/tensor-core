// module memory_arbiter #(
//   parameter BUS_SIZE = 32,      // General Bus Size
//   parameter MAT_BUS_SIZE = 64,      // Matrix Bus Size
// )(
//   input logic CLK, nRST
// );
  

// endmodule