// fust gets written do in dispatch on clock edge
// issue should read registers and issue to execute by the next clock edge
