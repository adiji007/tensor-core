//By            : Joe Nasti
//Last updated  : 11/17/2024 - reduced to 16 bit FP values for systolic array
//
//Module summary:
//    First step for addition operation in three-step pipline.
//    Shifts smaller fraction by difference in exponents
//
//Inputs:
//    floating_point1/2_in - single precision floating point values
//Outputs:
//    sign_shifted         - sign of the floating point that gets shifted
//    frac_shifted         - fraction of the floating point that gets shifted
//    sign_not_shifted     - sign of the floating point that does not get shifted
//    frac_not_shifted     - fraction of the floating point that does not get shifted
//    exp_max              - max exponent of the two given floating points

`timescale 1ns/1ps

module ADD_step1 (
    input  logic [15:0] floating_point1_in,
    input  logic [15:0] floating_point2_in,
    output logic sign_shifted,
    output logic [12:0] frac_shifted,
    output logic sign_not_shifted,
    output logic [12:0] frac_not_shifted,
    output logic [4:0] exp_max
);

    reg  [4:0]   unsigned_exp_diff;
    reg    cmp_out;

    // int_compare:
    // if exp1 >= exp2: cmp_out = 0
    // if exp2 > exp1: cmp_out = 1
    int_compare cmp_exponents (
        .exp1(floating_point1_in[14:10]),
        .exp2(floating_point2_in[14:10]),
        .u_diff(unsigned_exp_diff),
        .cmp_out(cmp_out)
    );
    
    // need to: right shift significand (fraction) of number with smaller exponent
    // Fraction format: {1'b1, fp_fraction[9:0], 2'b00}
    always_comb begin
        if(cmp_out == 1) begin
            frac_shifted = {1'b1, floating_point1_in[9:0], 2'b00} >> unsigned_exp_diff;
            sign_shifted = floating_point1_in[15];
            frac_not_shifted = {1'b1, floating_point2_in[9:0], 2'b00};
            sign_not_shifted = floating_point2_in[15];
            exp_max = floating_point2_in[14:10];
        end
        else begin
            frac_shifted = {1'b1, floating_point2_in[9:0], 2'b00} >> unsigned_exp_diff;
            sign_shifted = floating_point2_in[15];
            frac_not_shifted = {1'b1, floating_point1_in[9:0], 2'b00};
            sign_not_shifted = floating_point1_in[15];
            exp_max = floating_point1_in[14:10];
        end
    end

endmodule
