`timescale 1ns / 10ps
`include "isa_types.vh"
`include "datapath_types.vh"

`include "fetch_branch_if.vh"
`include "fetch_if.vh"
`include "fu_branch_predictor_if.vh"
`include "fu_branch_if.vh"

import isa_pkg::*;

module fetch_branch_tb;

    parameter PERIOD = 2;
    logic CLK = 0, nRST;
    logic ihit = 1;

  // clock
    always #(PERIOD/2) CLK++;


    fetch_branch_if fbif();
    fetch_if fif();
    fu_branch_predictor_if fubpif();
    fu_branch_if fubif();

    test PROG (CLK, nRST, fbif);

    fetch_branch FB (.CLK(CLK), .nRST(nRST), .fbif(fbif));
    fetch FETCH (.CLK(CLK), .nRST(nRST), .ihit(ihit), .fif(fif));
    fu_branch_predictor FUBR (.CLK(CLK), .nRST(nRST), .fubpif(fubpif));
    fu_branch FUB (.CLK(CLK), .nRST(nRST), .fubif(fubif));
endmodule 

    program test (input logic CLK, 
                  output logic nRST, 
                  fetch_branch_if.fb fbif);

    parameter CLOCK_TIME = 10;
    initial begin

    nRST = 0;
    fbif.imemload = '0;
    fbif.flush = '0;
    fbif.stall = '0;
    fbif.dispatch_free = '0;
    fbif.branch = '0;
    fbif.branch_type = 2'b00;
    fbif.branch_gate_sel = 1'b0;
    fbif.reg_a = 32'd0;
    fbif.reg_b = 32'd0;
    fbif.current_pc = 32'd0;
    fbif.imm = 32'd0;
    fbif.predicted_outcome = '0;
    fbif.current_pc = '0;

    @(posedge CLK);
    nRST = 1;

    #(CLOCK_TIME * 80);
    
    $finish;
    end
    endprogram 
 
