//thisdoesnt work