

// rishi doing control

module control_unit ();

endmodule